.control
    set wr_singlescale
    option numdgt = 4
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vth]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vdsat]
    
    run
    wrdata sweep_nmos_lvt_outchar.dat
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vth]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vdsat]
    
    save @m.xm1.msky130_fd_pr__nfet_01v8[id]
    save @m.xm1.msky130_fd_pr__nfet_01v8[vth]
    save @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
    
    run
    wrdata sweep_nmos_outchar.dat
    + @m.xm1.msky130_fd_pr__nfet_01v8[id]
    + @m.xm1.msky130_fd_pr__nfet_01v8[vth]
    + @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
.endc
