** sch_path: /home/ttuser/work/tt08-analog-template/work/design/nmos.sch
**.subckt nmos
XM1 VDS VGS VSS VBS sky130_fd_pr__nfet_01v8 L={L} W={W} nf={F} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult={M} m={M}
vgs VGS VSS 0
V4 VBS VSS {vbs}
V7 VSS GND 0
V8 VDS VSS {vds}
XM2 VDS VGS VSS VBS sky130_fd_pr__nfet_01v8_lvt L={L} W={W} nf={F} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult={M} m={M}
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice




.include nmos_param.spice
.include nmos_ctrl.spice



**** end user architecture code
**.ends
.GLOBAL GND
.end
