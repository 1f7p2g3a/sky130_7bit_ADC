.param Ln = 0.5
.param Wn = 10
.param Fn = 1
.param Mn = 1
.param Lp = 0.5
.param Wp = 10
.param Fp = 1
.param Mp = 1
.dc vin 0 1.8 0.01
