.control
    set wr_singlescale
    option numdgt = 4
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vth]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vdsat]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gmbs]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gds]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cbb]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[csb]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cdb]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cgb]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[css]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[csd]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[csg]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cds]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cdd]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cdg]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cbs]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cbd]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cbg]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cgd]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cgs]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cgg]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[capbs]
    save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[capbd]
    
    run
    wrdata sweep_nmos_lvt.dat
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vth]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vdsat]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gmbs]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gds]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cbb]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[csb]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cdb]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cgb]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[css]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[csd]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[csg]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cds]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cdd]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cdg]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cbs]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cbd]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cbg]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cgd]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cgs]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cgg]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[capbs]
    + @m.xm2.msky130_fd_pr__nfet_01v8_lvt[capbd]
    
    save @m.xm1.msky130_fd_pr__nfet_01v8[id]
    save @m.xm1.msky130_fd_pr__nfet_01v8[vth]
    save @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
    save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
    save @m.xm1.msky130_fd_pr__nfet_01v8[gmbs]
    save @m.xm1.msky130_fd_pr__nfet_01v8[gds]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cbb]
    save @m.xm1.msky130_fd_pr__nfet_01v8[csb]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cdb]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cgb]
    save @m.xm1.msky130_fd_pr__nfet_01v8[css]
    save @m.xm1.msky130_fd_pr__nfet_01v8[csd]
    save @m.xm1.msky130_fd_pr__nfet_01v8[csg]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cds]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cdd]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cdg]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cbs]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cbd]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cbg]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cgd]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cgs]
    save @m.xm1.msky130_fd_pr__nfet_01v8[cgg]
    save @m.xm1.msky130_fd_pr__nfet_01v8[capbs]
    save @m.xm1.msky130_fd_pr__nfet_01v8[capbd]
    
    run
    wrdata sweep_nmos.dat
    + @m.xm1.msky130_fd_pr__nfet_01v8[id]
    + @m.xm1.msky130_fd_pr__nfet_01v8[vth]
    + @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
    + @m.xm1.msky130_fd_pr__nfet_01v8[gm]
    + @m.xm1.msky130_fd_pr__nfet_01v8[gmbs]
    + @m.xm1.msky130_fd_pr__nfet_01v8[gds]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cbb]
    + @m.xm1.msky130_fd_pr__nfet_01v8[csb]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cdb]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cgb]
    + @m.xm1.msky130_fd_pr__nfet_01v8[css]
    + @m.xm1.msky130_fd_pr__nfet_01v8[csd]
    + @m.xm1.msky130_fd_pr__nfet_01v8[csg]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cds]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cdd]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cdg]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cbs]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cbd]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cbg]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cgd]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cgs]
    + @m.xm1.msky130_fd_pr__nfet_01v8[cgg]
    + @m.xm1.msky130_fd_pr__nfet_01v8[capbs]
    + @m.xm1.msky130_fd_pr__nfet_01v8[capbd]
.endc
