.param Wpm = 2.0
.param Lnm = 0.15
.param Lpm = 0.15
.param Wnm = 0.42
.param Fnm = 1
.param Mnm = 1
.param Fpm = 1
.param Mpm = 1
.dc vin 0 1.8 0.01